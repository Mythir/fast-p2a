-- Licensed under the Apache License, Version 2.0 (the "License");
-- you may not use this file except in compliance with the License.
-- You may obtain a copy of the License at
--
--     http://www.apache.org/licenses/LICENSE-2.0
--
-- Unless required by applicable law or agreed to in writing, software
-- distributed under the License is distributed on an "AS IS" BASIS,
-- WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
-- See the License for the specific language governing permissions and
-- limitations under the License.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
-- Fletcher utils, for use of log2ceil function.
use work.UtilInt_pkg.all;

-- This is a testbench for the ShifterRecombiner. The ShifterRecombiner will shift the bus words in its pipeline with a constant amount and then 
-- recombine the split bus words into complete (aligned) bus words.
-- If the alignment of the bus words changes while the ShifterRecombiner is already processing data the pipeline contents will have to be invalidated.
-- If there were any bus words in the pipeline that should have been shifted with the new alignment than those bus words will have to be re-entered into the pipeline.
-- (The testbench takes care of this.)

-- Use ShifterRecombiner_gen.py to generate ROM's containing misaligned data.

entity ShifterRecombiner_tb is
end ShifterRecombiner_tb;

architecture tb of ShifterRecombiner_tb is
  constant BUS_DATA_WIDTH         : natural := 512;
  constant ELEMENT_WIDTH          : natural := 8;
  constant SHIFT_WIDTH            : natural := log2ceil(BUS_DATA_WIDTH/ELEMENT_WIDTH);
  constant NUM_SHIFT_STAGES       : natural := SHIFT_WIDTH;
  constant clk_period                : time := 10 ns;

  signal clk                      : std_logic;
  signal reset                    : std_logic;
  signal clear                    : std_logic;
  signal in_valid                 : std_logic;
  signal in_ready                 : std_logic;
  signal in_data                  : std_logic_vector(BUS_DATA_WIDTH-1 downto 0);
  signal out_valid                : std_logic;
  signal out_ready                : std_logic;
  signal out_data                 : std_logic_vector(BUS_DATA_WIDTH-1 downto 0);
  signal alignment                : std_logic_vector(SHIFT_WIDTH-1 downto 0);

  -- Signals for checking output
  signal consumed_word            : std_logic_vector(BUS_DATA_WIDTH-1 downto 0);
  signal num_consumed_words       : integer;

  -- Misaligned input of the ShifterRecombiner
  type mem1 is array (0 to 33) of std_logic_vector(511 downto 0);
  constant MisalignedBusWord_ROM : mem1 := (
    0 => x"00000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
    1 => x"11111111222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222",
    2 => x"22222222333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333",
    3 => x"33333333444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444",
    4 => x"44444444555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555",
    5 => x"55555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555566",
    6 => x"66666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666677",
    7 => x"77777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777788",
    8 => x"88888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888899",
    9 => x"99999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999900",
    10 => x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011",
    11 => x"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111122",
    12 => x"22222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222233",
    13 => x"33333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333344",
    14 => x"44444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444455",
    15 => x"55555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555566",
    16 => x"77777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777",
    17 => x"88888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888",
    18 => x"99999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999",
    19 => x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
    20 => x"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
    21 => x"22222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222",
    22 => x"22222222222222222222222222222222222222222222222222222222222233333333333333333333333333333333333333333333333333333333333333333333",
    23 => x"33333333333333333333333333333333333333333333333333333333333344444444444444444444444444444444444444444444444444444444444444444444",
    24 => x"55555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555",
    25 => x"66666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666",
    26 => x"77777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777",
    27 => x"88888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888",
    28 => x"88888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888999999999999999999",
    29 => x"99999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999000000000000000000",
    30 => x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111",
    31 => x"22222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222",
    32 => x"33333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333",
    33 => x"44444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444"
  );
  
  --Alignment of all bus words in MisalignedBusWord_ROM
  type mem2 is array (0 to 33) of integer;
  constant Alignment_ROM : mem2 := (
    0 => 4,
    1 => 4,
    2 => 4,
    3 => 4,
    4 => 4,
    5 => 63,
    6 => 63,
    7 => 63,
    8 => 63,
    9 => 63,
    10 => 63,
    11 => 63,
    12 => 63,
    13 => 63,
    14 => 63,
    15 => 63,
    16 => 0,
    17 => 0,
    18 => 0,
    19 => 0,
    20 => 0,
    21 => 0,
    22 => 30,
    23 => 30,
    24 => 0,
    25 => 0,
    26 => 0,
    27 => 0,
    28 => 55,
    29 => 55,
    30 => 55,
    31 => 0,
    32 => 0,
    33 => 0
  );
  
  --List of aligned bus words we expect the ShifterRecombiner to produce
  type mem3 is array (0 to 29) of std_logic_vector(511 downto 0);
  constant AlignedBusWord_ROM : mem3 := (
    0 => x"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
    1 => x"22222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222",
    2 => x"33333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333",
    3 => x"44444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444",
    4 => x"66666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666",
    5 => x"77777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777",
    6 => x"88888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888",
    7 => x"99999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999",
    8 => x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
    9 => x"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
    10 => x"22222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222",
    11 => x"33333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333",
    12 => x"44444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444",
    13 => x"55555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555",
    14 => x"77777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777",
    15 => x"88888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888",
    16 => x"99999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999",
    17 => x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
    18 => x"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
    19 => x"22222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222",
    20 => x"33333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333",
    21 => x"55555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555",
    22 => x"66666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666",
    23 => x"77777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777",
    24 => x"88888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888",
    25 => x"99999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999",
    26 => x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
    27 => x"22222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222",
    28 => x"33333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333",
    29 => x"44444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444"
  );
  
  --Original alignment of all bus words in AlignedBusWord_ROM
  type mem4 is array (0 to 29) of integer;
  constant Alignment2_ROM : mem4 := (
    0 => 4,
    1 => 4,
    2 => 4,
    3 => 4,
    4 => 63,
    5 => 63,
    6 => 63,
    7 => 63,
    8 => 63,
    9 => 63,
    10 => 63,
    11 => 63,
    12 => 63,
    13 => 63,
    14 => 0,
    15 => 0,
    16 => 0,
    17 => 0,
    18 => 0,
    19 => 0,
    20 => 30,
    21 => 0,
    22 => 0,
    23 => 0,
    24 => 0,
    25 => 55,
    26 => 55,
    27 => 0,
    28 => 0,
    29 => 0
  );

begin
  dut: entity work.ShifterRecombiner
  generic map(
    BUS_DATA_WIDTH              => BUS_DATA_WIDTH,
    SHIFT_WIDTH                 => SHIFT_WIDTH,
    ELEMENT_WIDTH               => ELEMENT_WIDTH,
    NUM_SHIFT_STAGES            => NUM_SHIFT_STAGES
  )
  port map(
    clk                         => clk,
    reset                       => reset,
    clear                       => clear,
    in_valid                    => in_valid,
    in_ready                    => in_ready,
    in_data                     => in_data,
    out_valid                   => out_valid,
    out_ready                   => out_ready,
    out_data                    => out_data,
    alignment                   => alignment
  );

  -- This process is responsible for data input into the ShifterRecombiner
  upstream_p : process
    -- Current index for input data
    variable i : integer := 0;

    -- Amount of times we had to realign
    variable realignments : integer := 0;
  begin
    in_valid <= '0';
    loop
      wait until rising_edge(clk);
      exit when reset = '0';
    end loop;

    -- Starting alignment
    alignment <= std_logic_vector(to_unsigned(Alignment_ROM(i), alignment'length));

    loop
      -- Downstream signals an alignment change with the clear signal.
      if clear = '1' then
        -- Alignment change        

        -- A little bit gross: when alignment is zero there is an extra valid bus word. Therefore, when the previous alignment was 0, we decrement
        -- the amount of realignments to ensure the input data starts from the correct index again.
        if to_integer(unsigned(alignment)) = 0 then
          realignments := realignments - 1;
        end if;

        alignment <= std_logic_vector(to_unsigned(Alignment_ROM(num_consumed_words + realignments + 1), alignment'length));
        -- The testbench simulates the case where the hardware around the ShifterRecombiner knows in what bus word the alignment changes
        i := num_consumed_words + realignments + 1;
        realignments := realignments + 1;
      end if;

      -- Avoid reading data out of the range of the MisalignedBusWord_ROM
      if i < MisalignedBusWord_ROM'length then
        in_valid <= '1';
        in_data <= MisalignedBusWord_ROM(i);
  
        loop
          wait until rising_edge(clk);
          exit when in_ready = '1';
        end loop;
      else
        wait until rising_edge(clk);
      end if;

      in_valid <= '0';

      i := i+1;
    end loop;
    wait;
  end process;

  -- This process is responsible for consuming the ShifterRecombiner output data and checking it's correctness.
  downstream_p : process
    -- Current index in the ROM with expected results
    variable j : integer := 0;
  begin
    num_consumed_words <= 0;
    clear <= '0';
    out_ready <= '0';
    loop
      wait until rising_edge(clk);
      exit when reset = '0';
    end loop;

    loop
      clear <= '0';

      out_ready <= '1';

      loop
        wait until rising_edge(clk);
        exit when out_valid = '1';
      end loop;

      consumed_word <= out_data;
      num_consumed_words <= num_consumed_words + 1;
      out_ready <= '0';

      -- Automatic output check
      assert out_data = AlignedBusWord_ROM(j)
        report "Unexpected output at aligned bus word " & integer'image(j);

      if j+1 < Alignment2_ROM'length then
        if Alignment2_ROM(j+1) /= Alignment2_ROM(j) then
          -- Signal alignment change
          clear <= '1';
          wait until rising_edge(clk);
        end if;
      end if;

      j := j+1;

      -- Exit this loop when all expected words have been read
      exit when j = AlignedBusWord_ROM'length;
    end loop;
    report "Simulation completed successfully";
    wait;
  end process;

  clk_p : process
  begin
    clk <= '0';
    wait for clk_period/2;
    clk <= '1';
    wait for clk_period/2;
  end process;

  reset_p : process is
  begin
    reset <= '1';
    wait for 20 ns;
    wait until rising_edge(clk);
    reset <= '0';
    wait;
  end process;
end architecture;

-- Copyright 2018 Delft University of Technology
--
-- Licensed under the Apache License, Version 2.0 (the "License");
-- you may not use this file except in compliance with the License.
-- You may obtain a copy of the License at
--
--     http://www.apache.org/licenses/LICENSE-2.0
--
-- Unless required by applicable law or agreed to in writing, software
-- distributed under the License is distributed on an "AS IS" BASIS,
-- WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
-- See the License for the specific language governing permissions and
-- limitations under the License.

library std;
use std.textio.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_textio.all;
use ieee.math_real.all;

library work;
-- Fletcher utils, for use of log2ceil function.
use work.UtilInt_pkg.all;

-- This testbench takes input generated by the V2MetadataInterpreter_gen.py and streams it into the MetadataInterpreter.
-- Using the correct output files from the Python script this testbench then verifies that the MetadataInterpreter functions
-- correctly.
-- This testbench also sometimes stops the input stream for a random amount of cycles to check the MetadataInterpreter under
-- non-continuous input stream conditions.

entity V2MetadataInterpreter_tb is
end V2MetadataInterpreter_tb;

architecture tb of V2MetadataInterpreter_tb is
  constant clk_period                : time    := 10 ns;
  constant BUS_DATA_WIDTH            : natural := 512;
  constant CYCLE_COUNT_WIDTH         : natural := 8;

  -- Probability of an interruption in the input stream
  constant stream_stop_p        : real    := 0.20;
  -- Max amount of stopped cycles in case of an interruption
  constant max_stopped_cycles   : real    := 75.0;

  signal clk                         : std_logic;
  signal hw_reset                    : std_logic;
  signal in_valid                    : std_logic;
  signal in_ready                    : std_logic;
  signal in_data                     : std_logic_vector(BUS_DATA_WIDTH-1 downto 0);
  signal da_valid                    : std_logic;
  signal da_ready                    : std_logic;
  signal da_bytes_consumed           : std_logic_vector(log2ceil(BUS_DATA_WIDTH/8) downto 0);
  signal rl_byte_length              : std_logic_vector(31 downto 0);
  signal dl_byte_length              : std_logic_vector(31 downto 0);
  signal dc_uncomp_size              : std_logic_vector(31 downto 0);
  signal dc_comp_size                : std_logic_vector(31 downto 0);
  signal dd_num_values               : std_logic_vector(31 downto 0);

begin
  dut : entity work.V2MetadataInterpreter
  generic map(
    BUS_DATA_WIDTH => BUS_DATA_WIDTH
  )
  port map(
    clk                 => clk,
    hw_reset            => hw_reset,
    in_valid            => in_valid,
    in_ready            => in_ready,
    in_data             => in_data,
    da_valid            => da_valid,
    da_ready            => da_ready,
    da_bytes_consumed   => da_bytes_consumed,
    rl_byte_length      => rl_byte_length,
    dl_byte_length      => dl_byte_length,
    dc_uncomp_size      => dc_uncomp_size,
    dc_comp_size        => dc_comp_size,
    dd_num_values       => dd_num_values
  );

  upstream_p: process is
    file input_data             : text;

    variable input_line         : line;
    variable bus_word           : std_logic_vector(BUS_DATA_WIDTH-1 downto 0);

    variable seed1              : positive := 1337;
    variable seed2              : positive := 4242;

    variable stream_stop        : real;
    variable num_stopped_cycles : real;
  begin
    file_open(input_data, "./test/thrift/V2MDI_input.hex", read_mode);
    in_valid <= '0';

    loop
      wait until rising_edge(clk);
      exit when hw_reset = '0';
    end loop;

    while not endfile(input_data) loop
      readline(input_data, input_line);
      hread(input_line, bus_word);

      in_valid <= '1';
      in_data <= bus_word;
  
      loop
        wait until rising_edge(clk);
        exit when in_ready = '1';
      end loop;
  
      in_valid <= '0';

      -- Delay for a random amount of clock cycles to simulate a non-continuous stream
      uniform(seed1, seed2, stream_stop);
      if stream_stop < stream_stop_p then
        uniform(seed1, seed2, num_stopped_cycles);
        for i in 0 to integer(floor(num_stopped_cycles*max_stopped_cycles)) loop
          wait until rising_edge(clk);
        end loop;
      end if;
    end loop;

    report "All metadata input has been processed";

    wait;
  end process;

  downstream_p: process is
    file output_data             : text;

    variable output_line         : line;
    variable space               : character;

    variable uncomp_size         : std_logic_vector(31 downto 0);
    variable comp_size           : std_logic_vector(31 downto 0);
    variable num_val             : std_logic_vector(31 downto 0);
    variable def_lvl             : std_logic_vector(31 downto 0);
    variable rep_lvl             : std_logic_vector(31 downto 0);
  begin
    file_open(output_data, "./test/thrift/V2MDI_output.hex", read_mode);
    da_ready <= '0';

    loop
      wait until rising_edge(clk);
      exit when hw_reset = '0';
    end loop;

    while not endfile(output_data) loop
      readline(output_data, output_line);
      hread(output_line, uncomp_size);
      read(output_line, space);
      hread(output_line, comp_size);
      read(output_line, space);
      hread(output_line, num_val);
      read(output_line, space);
      hread(output_line, def_lvl);
      read(output_line, space);
      hread(output_line, rep_lvl);

      da_ready <= '1';

      loop
        wait until rising_edge(clk);
        exit when da_valid = '1';
      end loop;

      assert uncomp_size = dc_uncomp_size
        report "uncomp_size = " & integer'image(to_integer(unsigned(dc_uncomp_size))) & ", should be " & integer'image(to_integer(unsigned(uncomp_size))) severity failure;
      assert comp_size = dc_comp_size
        report "comp_size = " & integer'image(to_integer(unsigned(dc_comp_size))) & ", should be " & integer'image(to_integer(unsigned(comp_size))) severity failure;
      assert num_val = dd_num_values
        report "num_val = " & integer'image(to_integer(unsigned(dd_num_values))) & ", should be " & integer'image(to_integer(unsigned(num_val))) severity failure;
      assert def_lvl = dl_byte_length
        report "dl byte length = " & integer'image(to_integer(unsigned(dl_byte_length))) & ", should be " & integer'image(to_integer(unsigned(def_lvl))) severity failure;
      assert rep_lvl = rl_byte_length
        report "rl byte length = " & integer'image(to_integer(unsigned(rl_byte_length))) & ", should be " & integer'image(to_integer(unsigned(rep_lvl))) severity failure;

      da_ready <= '0';
    end loop;

    report "All metadata output has been processed";

    wait;
  end process;

  clk_p :process
  begin
    clk <= '0';
    wait for clk_period/2;
    clk <= '1';
    wait for clk_period/2;
  end process;

  reset_p: process is
  begin
    hw_reset <= '1';
    wait for 20 ns;
    wait until rising_edge(clk);
    hw_reset <= '0';
    wait;
  end process;
end architecture;
